
module nes_test_controller ();



endmodule